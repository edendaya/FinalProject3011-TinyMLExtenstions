// Verilog test fixture created from schematic E:\adlx\D4\monitor\monitor.sch - Mon Nov 25 14:45:29 2024

`timescale 1ns / 1ps

module monitor_monitor_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   monitor UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:08:25 11/18/2024 
// Design Name: 
// Module Name:    ID_NUM 
// Project Name: 
// Target Devices: 

// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ID_NUM(
		output [7:0] ID
    );
	 assign ID = 8'hD4;
	 

endmodule
